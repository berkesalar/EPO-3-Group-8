library ieee;
use ieee.std_logic_1164.all;

entity level_lut is
    port (
        addr    : in std_logic_vector(11 downto 0);
        blk_data: out std_logic_vector(3 downto 0)
    );
end entity level_lut;


architecture lut of level_lut is

begin

    -- Sprite (2 bits) & collision data (2 bits) in each 16x21 screen:
    -- Sprite: 00-- = air, 01-- = brick, 10-- = block;
    -- Collision: --00 = no collision, --01 = collision, --10 = death, --11 = win
    with addr select blk_data <=
        -- all blocks except 'air' in screen 0 are below
        "1001" when "000000000000",  -- brick
        "1001" when "000011010010",  -- brick
        "1001" when "000110100100",  -- brick
        "1001" when "001001110110",  -- brick
        "1001" when "001101001000",  -- brick
        "1001" when "010000011010",  -- brick
        "1001" when "010011101100",  -- brick
        "1001" when "010110111110",  -- brick
        "1001" when "011010010000",  -- brick
        "1001" when "011101100010",  -- brick
        "1001" when "100000110100",  -- brick
        "1001" when "100100000110",  -- brick
        "1001" when "100111011000",  -- brick
        "0101" when "101010101010",  -- block
        "0101" when "101101111100",  -- block
        "0010" when "110001001110",  -- death
        "0101" when "101010101011",  -- block
        "0101" when "101101111101",  -- block
        "0010" when "110001001111",  -- death
        "0101" when "101010101100",  -- block
        "0101" when "101101111110",  -- block
        "0010" when "110001010000",  -- death
        "0101" when "101010101101",  -- block
        "0101" when "101101111111",  -- block
        "0010" when "110001010001",  -- death
        "0101" when "101010101110",  -- block
        "0101" when "101110000000",  -- block
        "0010" when "110001010010",  -- death
        "0101" when "101010101111",  -- block
        "0101" when "101110000001",  -- block
        "0010" when "110001010011",  -- death
        "0101" when "101010110000",  -- block
        "0101" when "101110000010",  -- block
        "0010" when "110001010100",  -- death
        "0101" when "101010110001",  -- block
        "0101" when "101110000011",  -- block
        "0010" when "110001010101",  -- death
        "0101" when "101010110010",  -- block
        "0101" when "101110000100",  -- block
        "0010" when "110001010110",  -- death
        "0101" when "101010110011",  -- block
        "0101" when "101110000101",  -- block
        "0010" when "110001010111",  -- death
        "0101" when "101010110100",  -- block
        "0101" when "101110000110",  -- block
        "0010" when "110001011000",  -- death
        "0101" when "101010110101",  -- block
        "0101" when "101110000111",  -- block
        "0010" when "110001011001",  -- death
        "0101" when "101010110110",  -- block
        "0101" when "101110001000",  -- block
        "0010" when "110001011010",  -- death
        "0101" when "101010110111",  -- block
        "0101" when "101110001001",  -- block
        "0010" when "110001011011",  -- death
        "0101" when "101010111000",  -- block
        "0101" when "101110001010",  -- block
        "0010" when "110001011100",  -- death
        "0101" when "101010111001",  -- block
        "0101" when "101110001011",  -- block
        "0010" when "110001011101",  -- death
        "0101" when "101010111010",  -- block
        "0101" when "101110001100",  -- block
        "0010" when "110001011110",  -- death
        "1001" when "011101110011",  -- brick
        "0101" when "101010111011",  -- block
        "0101" when "101110001101",  -- block
        "0010" when "110001011111",  -- death
        "0101" when "101010111100",  -- block
        "0101" when "101110001110",  -- block
        "0010" when "110001100000",  -- death
        "0101" when "101010111101",  -- block
        "0101" when "101110001111",  -- block
        "0010" when "110001100001",  -- death
        "0101" when "101010111110",  -- block
        "0101" when "101110010000",  -- block
        "0010" when "110001100010",  -- death
        -- all blocks except 'air' in screen 1 are below
        "1001" when "011101110111",  -- brick
        "0101" when "101010111111",  -- block
        "0101" when "101110010001",  -- block
        "0010" when "110001100011",  -- death
        "0101" when "011101111000",  -- block
        "0101" when "101011000000",  -- block
        "0101" when "101110010010",  -- block
        "0010" when "110001100100",  -- death
        "0101" when "010000110001",  -- block
        "1001" when "011101111001",  -- brick
        "0101" when "101011000001",  -- block
        "0101" when "101110010011",  -- block
        "0010" when "110001100101",  -- death
        "0101" when "011101111010",  -- block
        "0101" when "101011000010",  -- block
        "0101" when "101110010100",  -- block
        "0010" when "110001100110",  -- death
        "1001" when "011101111011",  -- brick
        "0101" when "101011000011",  -- block
        "0101" when "101110010101",  -- block
        "0010" when "110001100111",  -- death
        "0101" when "101011000100",  -- block
        "0101" when "101110010110",  -- block
        "0010" when "110001101000",  -- death
        "0101" when "101011000101",  -- block
        "0101" when "101110010111",  -- block
        "0010" when "110001101001",  -- death
        "0101" when "101011000110",  -- block
        "0101" when "101110011000",  -- block
        "0010" when "110001101010",  -- death
        "1001" when "100100100011",  -- brick
        "1001" when "100111110101",  -- brick
        "0101" when "101011000111",  -- block
        "0101" when "101110011001",  -- block
        "0010" when "110001101011",  -- death
        "1001" when "100100100100",  -- brick
        "1001" when "100111110110",  -- brick
        "0101" when "101011001000",  -- block
        "0101" when "101110011010",  -- block
        "0010" when "110001101100",  -- death
        "0101" when "101011001001",  -- block
        "0101" when "101110011011",  -- block
        "0010" when "110001101101",  -- death
        "0101" when "101011001010",  -- block
        "0101" when "101110011100",  -- block
        "0010" when "110001101110",  -- death
        "0101" when "101011001011",  -- block
        "0101" when "101110011101",  -- block
        "0010" when "110001101111",  -- death
        "0101" when "101011001100",  -- block
        "0101" when "101110011110",  -- block
        "0010" when "110001110000",  -- death
        "0101" when "101011001101",  -- block
        "0101" when "101110011111",  -- block
        "0010" when "110001110001",  -- death
        "0101" when "101011001110",  -- block
        "0101" when "101110100000",  -- block
        "0010" when "110001110010",  -- death
        "0101" when "101011001111",  -- block
        "0101" when "101110100001",  -- block
        "0010" when "110001110011",  -- death
        "1001" when "100001011010",  -- brick
        "0101" when "101011010000",  -- block
        "0101" when "101110100010",  -- block
        "0010" when "110001110100",  -- death
        "1001" when "100001011011",  -- brick
        "1001" when "100100101101",  -- brick
        "1001" when "100111111111",  -- brick
        "0101" when "101011010001",  -- block
        "0101" when "101110100011",  -- block
        "0010" when "110001110101",  -- death
        "1001" when "100001011100",  -- brick
        "1001" when "100100101110",  -- brick
        "1001" when "101000000000",  -- brick
        "0101" when "101011010010",  -- block
        "0101" when "101110100100",  -- block
        "0010" when "110001110110",  -- death
        "1001" when "100001011101",  -- brick
        "0101" when "101011010011",  -- block
        "0101" when "101110100101",  -- block
        "0010" when "110001110111",  -- death
        -- all blocks except 'air' in screen 2 are below
        "0101" when "101011010100",  -- block
        "0101" when "101110100110",  -- block
        "0010" when "110001111000",  -- death
        "0101" when "101011010101",  -- block
        "0101" when "101110100111",  -- block
        "0010" when "110001111001",  -- death
        "0101" when "101011010110",  -- block
        "0101" when "101110101000",  -- block
        "0010" when "110001111010",  -- death
        "0101" when "101011010111",  -- block
        "0101" when "101110101001",  -- block
        "0010" when "110001111011",  -- death
        "1001" when "011110010000",  -- brick
        "0101" when "101011011000",  -- block
        "0101" when "101110101010",  -- block
        "0010" when "110001111100",  -- death
        "1001" when "011110010001",  -- brick
        "1001" when "100001100011",  -- brick
        "1001" when "100100110101",  -- brick
        "1001" when "101000000111",  -- brick
        "0101" when "101011011001",  -- block
        "0101" when "101110101011",  -- block
        "0010" when "110001111101",  -- death
        "1001" when "011110010010",  -- brick
        "1001" when "100001100100",  -- brick
        "1001" when "100100110110",  -- brick
        "1001" when "101000001000",  -- brick
        "0101" when "101011011010",  -- block
        "0101" when "101110101100",  -- block
        "0010" when "110001111110",  -- death
        "1001" when "011110010011",  -- brick
        "0101" when "101011011011",  -- block
        "0101" when "101110101101",  -- block
        "0010" when "110001111111",  -- death
        "0101" when "101011011100",  -- block
        "0101" when "101110101110",  -- block
        "0010" when "110010000000",  -- death
        "0101" when "101011011101",  -- block
        "0101" when "101110101111",  -- block
        "0010" when "110010000001",  -- death
        "0101" when "101011011110",  -- block
        "0101" when "101110110000",  -- block
        "0010" when "110010000010",  -- death
        "0101" when "101011011111",  -- block
        "0101" when "101110110001",  -- block
        "0010" when "110010000011",  -- death
        "0101" when "101011100000",  -- block
        "0101" when "101110110010",  -- block
        "0010" when "110010000100",  -- death
        "0101" when "101011100001",  -- block
        "0101" when "101110110011",  -- block
        "0010" when "110010000101",  -- death
        "0101" when "101011100010",  -- block
        "0101" when "101110110100",  -- block
        "0010" when "110010000110",  -- death
        "1001" when "011110011011",  -- brick
        "0101" when "101011100011",  -- block
        "0101" when "101110110101",  -- block
        "0010" when "110010000111",  -- death
        "1001" when "011110011100",  -- brick
        "1001" when "100001101110",  -- brick
        "1001" when "100101000000",  -- brick
        "1001" when "101000010010",  -- brick
        "0101" when "101011100100",  -- block
        "0101" when "101110110110",  -- block
        "0010" when "110010001000",  -- death
        "1001" when "011110011101",  -- brick
        "1001" when "100001101111",  -- brick
        "1001" when "100101000001",  -- brick
        "1001" when "101000010011",  -- brick
        "0101" when "101011100101",  -- block
        "0101" when "101110110111",  -- block
        "0010" when "110010001001",  -- death
        "1001" when "011110011110",  -- brick
        "0101" when "101011100110",  -- block
        "0101" when "101110111000",  -- block
        "0010" when "110010001010",  -- death
        "0101" when "101011100111",  -- block
        "0101" when "101110111001",  -- block
        "0010" when "110010001011",  -- death
        "0101" when "101011101000",  -- block
        "0101" when "101110111010",  -- block
        "0010" when "110010001100",  -- death
        -- all blocks except 'air' in screen 3 are below
        "0101" when "101011101001",  -- block
        "0101" when "101110111011",  -- block
        "0010" when "110010001101",  -- death
        "0101" when "101011101010",  -- block
        "0101" when "101110111100",  -- block
        "0010" when "110010001110",  -- death
        "0101" when "101011101011",  -- block
        "0101" when "101110111101",  -- block
        "0010" when "110010001111",  -- death
        "0101" when "101011101100",  -- block
        "0101" when "101110111110",  -- block
        "0010" when "110010010000",  -- death
        "0101" when "101011101101",  -- block
        "0101" when "101110111111",  -- block
        "0010" when "110010010001",  -- death
        "0101" when "101011101110",  -- block
        "0101" when "101111000000",  -- block
        "0010" when "110010010010",  -- death
        "0101" when "101011101111",  -- block
        "0101" when "101111000001",  -- block
        "0010" when "110010010011",  -- death
        "0010" when "110010010100",  -- death
        "0010" when "110010010101",  -- death
        "0101" when "101011110010",  -- block
        "0101" when "101111000100",  -- block
        "0010" when "110010010110",  -- death
        "0101" when "101011110011",  -- block
        "0101" when "101111000101",  -- block
        "0010" when "110010010111",  -- death
        "0101" when "101011110100",  -- block
        "0101" when "101111000110",  -- block
        "0010" when "110010011000",  -- death
        "0101" when "101011110101",  -- block
        "0101" when "101111000111",  -- block
        "0010" when "110010011001",  -- death
        "0101" when "101011110110",  -- block
        "0101" when "101111001000",  -- block
        "0010" when "110010011010",  -- death
        "0101" when "101011110111",  -- block
        "0101" when "101111001001",  -- block
        "0010" when "110010011011",  -- death
        "1001" when "011110110000",  -- brick
        "0101" when "101011111000",  -- block
        "0101" when "101111001010",  -- block
        "0010" when "110010011100",  -- death
        "0101" when "011110110001",  -- block
        "0101" when "101011111001",  -- block
        "0101" when "101111001011",  -- block
        "0010" when "110010011101",  -- death
        "1001" when "011110110010",  -- brick
        "0101" when "101011111010",  -- block
        "0101" when "101111001100",  -- block
        "0010" when "110010011110",  -- death
        "1001" when "010001101011",  -- brick
        "0101" when "101011111011",  -- block
        "0101" when "101111001101",  -- block
        "0010" when "110010011111",  -- death
        "1001" when "010001101100",  -- brick
        "0101" when "101011111100",  -- block
        "0101" when "101111001110",  -- block
        "0010" when "110010100000",  -- death
        "1001" when "010001101101",  -- brick
        "0101" when "101011111101",  -- block
        "0101" when "101111001111",  -- block
        "0010" when "110010100001",  -- death
        -- all blocks except 'air' in screen 4 are below
        "1001" when "010001101110",  -- brick
        "0101" when "101011111110",  -- block
        "0101" when "101111010000",  -- block
        "0010" when "110010100010",  -- death
        "1001" when "010001101111",  -- brick
        "0101" when "101011111111",  -- block
        "0101" when "101111010001",  -- block
        "0010" when "110010100011",  -- death
        "1001" when "010001110000",  -- brick
        "0101" when "101100000000",  -- block
        "0101" when "101111010010",  -- block
        "0010" when "110010100100",  -- death
        "1001" when "010001110001",  -- brick
        "0010" when "110010100101",  -- death
        "1001" when "010001110010",  -- brick
        "0010" when "110010100110",  -- death
        "0010" when "110010100111",  -- death
        "0101" when "101100000100",  -- block
        "0101" when "101111010110",  -- block
        "0010" when "110010101000",  -- death
        "0101" when "101100000101",  -- block
        "0101" when "101111010111",  -- block
        "0010" when "110010101001",  -- death
        "1001" when "010001110110",  -- brick
        "0101" when "101100000110",  -- block
        "0101" when "101111011000",  -- block
        "0010" when "110010101010",  -- death
        "1001" when "010001110111",  -- brick
        "0101" when "101100000111",  -- block
        "0101" when "101111011001",  -- block
        "0010" when "110010101011",  -- death
        "0101" when "010001111000",  -- block
        "1001" when "011111000000",  -- brick
        "0101" when "101100001000",  -- block
        "0101" when "101111011010",  -- block
        "0010" when "110010101100",  -- death
        "0101" when "101100001001",  -- block
        "0101" when "101111011011",  -- block
        "0010" when "110010101101",  -- death
        "0101" when "101100001010",  -- block
        "0101" when "101111011100",  -- block
        "0010" when "110010101110",  -- death
        "0101" when "101100001011",  -- block
        "0101" when "101111011101",  -- block
        "0010" when "110010101111",  -- death
        "0101" when "101100001100",  -- block
        "0101" when "101111011110",  -- block
        "0010" when "110010110000",  -- death
        "0101" when "101100001101",  -- block
        "0101" when "101111011111",  -- block
        "0010" when "110010110001",  -- death
        "1001" when "011111000110",  -- brick
        "0101" when "101100001110",  -- block
        "0101" when "101111100000",  -- block
        "0010" when "110010110010",  -- death
        "1001" when "011111000111",  -- brick
        "0101" when "101100001111",  -- block
        "0101" when "101111100001",  -- block
        "0010" when "110010110011",  -- death
        "0101" when "101100010000",  -- block
        "0101" when "101111100010",  -- block
        "0010" when "110010110100",  -- death
        "0101" when "101100010001",  -- block
        "0101" when "101111100011",  -- block
        "0010" when "110010110101",  -- death
        "0101" when "101100010010",  -- block
        "0101" when "101111100100",  -- block
        "0010" when "110010110110",  -- death
        -- all blocks except 'air' in screen 5 are below
        "0101" when "011111001011",  -- block
        "0101" when "101100010011",  -- block
        "0101" when "101111100101",  -- block
        "0010" when "110010110111",  -- death
        "0101" when "101100010100",  -- block
        "0101" when "101111100110",  -- block
        "0010" when "110010111000",  -- death
        "0101" when "101100010101",  -- block
        "0101" when "101111100111",  -- block
        "0010" when "110010111001",  -- death
        "0101" when "010010000110",  -- block
        "0101" when "011111001110",  -- block
        "0101" when "101100010110",  -- block
        "0101" when "101111101000",  -- block
        "0010" when "110010111010",  -- death
        "0101" when "101100010111",  -- block
        "0101" when "101111101001",  -- block
        "0010" when "110010111011",  -- death
        "0101" when "101100011000",  -- block
        "0101" when "101111101010",  -- block
        "0010" when "110010111100",  -- death
        "0101" when "011111010001",  -- block
        "0101" when "101100011001",  -- block
        "0101" when "101111101011",  -- block
        "0010" when "110010111101",  -- death
        "0101" when "101100011010",  -- block
        "0101" when "101111101100",  -- block
        "0010" when "110010111110",  -- death
        "0101" when "101100011011",  -- block
        "0101" when "101111101101",  -- block
        "0010" when "110010111111",  -- death
        "0101" when "101100011100",  -- block
        "0101" when "101111101110",  -- block
        "0010" when "110011000000",  -- death
        "0101" when "101100011101",  -- block
        "0101" when "101111101111",  -- block
        "0010" when "110011000001",  -- death
        "0101" when "101100011110",  -- block
        "0101" when "101111110000",  -- block
        "0010" when "110011000010",  -- death
        "1001" when "011111010111",  -- brick
        "0101" when "101100011111",  -- block
        "0101" when "101111110001",  -- block
        "0010" when "110011000011",  -- death
        "0101" when "101100100000",  -- block
        "0101" when "101111110010",  -- block
        "0010" when "110011000100",  -- death
        "0101" when "101100100001",  -- block
        "0101" when "101111110011",  -- block
        "0010" when "110011000101",  -- death
        "1001" when "010010010010",  -- brick
        "0101" when "101100100010",  -- block
        "0101" when "101111110100",  -- block
        "0010" when "110011000110",  -- death
        "1001" when "010010010011",  -- brick
        "0101" when "101100100011",  -- block
        "0101" when "101111110101",  -- block
        "0010" when "110011000111",  -- death
        "1001" when "010010010100",  -- brick
        "0101" when "101100100100",  -- block
        "0101" when "101111110110",  -- block
        "0010" when "110011001000",  -- death
        "0101" when "101100100101",  -- block
        "0101" when "101111110111",  -- block
        "0010" when "110011001001",  -- death
        "0101" when "101100100110",  -- block
        "0101" when "101111111000",  -- block
        "0010" when "110011001010",  -- death
        "0101" when "101100100111",  -- block
        "0101" when "101111111001",  -- block
        "0010" when "110011001011",  -- death
        -- all blocks except 'air' in screen 6 are below
        "0101" when "101100101000",  -- block
        "0101" when "101111111010",  -- block
        "0010" when "110011001100",  -- death
        "1001" when "010010011001",  -- brick
        "0101" when "101100101001",  -- block
        "0101" when "101111111011",  -- block
        "0010" when "110011001101",  -- death
        "0101" when "010010011010",  -- block
        "1001" when "011111100010",  -- brick
        "0101" when "101100101010",  -- block
        "0101" when "101111111100",  -- block
        "0010" when "110011001110",  -- death
        "0101" when "010010011011",  -- block
        "1001" when "011111100011",  -- brick
        "0101" when "101100101011",  -- block
        "0101" when "101111111101",  -- block
        "0010" when "110011001111",  -- death
        "1001" when "010010011100",  -- brick
        "0101" when "101100101100",  -- block
        "0101" when "101111111110",  -- block
        "0010" when "110011010000",  -- death
        "0101" when "101100101101",  -- block
        "0101" when "101111111111",  -- block
        "0010" when "110011010001",  -- death
        "0101" when "101100101110",  -- block
        "0101" when "110000000000",  -- block
        "0010" when "110011010010",  -- death
        "1001" when "101001011101",  -- brick
        "0101" when "101100101111",  -- block
        "0101" when "110000000001",  -- block
        "0010" when "110011010011",  -- death
        "1001" when "100110001100",  -- brick
        "1001" when "101001011110",  -- brick
        "0101" when "101100110000",  -- block
        "0101" when "110000000010",  -- block
        "0010" when "110011010100",  -- death
        "1001" when "100010111011",  -- brick
        "1001" when "100110001101",  -- brick
        "1001" when "101001011111",  -- brick
        "0101" when "101100110001",  -- block
        "0101" when "110000000011",  -- block
        "0010" when "110011010101",  -- death
        "1001" when "011111101010",  -- brick
        "1001" when "100010111100",  -- brick
        "1001" when "100110001110",  -- brick
        "1001" when "101001100000",  -- brick
        "0101" when "101100110010",  -- block
        "0101" when "110000000100",  -- block
        "0010" when "110011010110",  -- death
        "0101" when "101100110011",  -- block
        "0101" when "110000000101",  -- block
        "0010" when "110011010111",  -- death
        "0101" when "101100110100",  -- block
        "0101" when "110000000110",  -- block
        "0010" when "110011011000",  -- death
        "1001" when "011111101101",  -- brick
        "1001" when "100010111111",  -- brick
        "1001" when "100110010001",  -- brick
        "1001" when "101001100011",  -- brick
        "0101" when "101100110101",  -- block
        "0101" when "110000000111",  -- block
        "0010" when "110011011001",  -- death
        "1001" when "100011000000",  -- brick
        "1001" when "100110010010",  -- brick
        "1001" when "101001100100",  -- brick
        "0101" when "101100110110",  -- block
        "0101" when "110000001000",  -- block
        "0010" when "110011011010",  -- death
        "1001" when "100110010011",  -- brick
        "1001" when "101001100101",  -- brick
        "0101" when "101100110111",  -- block
        "0101" when "110000001001",  -- block
        "0010" when "110011011011",  -- death
        "1001" when "101001100110",  -- brick
        "0101" when "101100111000",  -- block
        "0101" when "110000001010",  -- block
        "0010" when "110011011100",  -- death
        "0101" when "101100111001",  -- block
        "0101" when "110000001011",  -- block
        "0010" when "110011011101",  -- death
        "0101" when "101100111010",  -- block
        "0101" when "110000001100",  -- block
        "0010" when "110011011110",  -- death
        "0101" when "101100111011",  -- block
        "0101" when "110000001101",  -- block
        "0010" when "110011011111",  -- death
        "0101" when "101100111100",  -- block
        "0101" when "110000001110",  -- block
        "0010" when "110011100000",  -- death
        -- all blocks except 'air' in screen 7 are below
        "1001" when "101001101011",  -- brick
        "0101" when "101100111101",  -- block
        "0101" when "110000001111",  -- block
        "0010" when "110011100001",  -- death
        "1001" when "100110011010",  -- brick
        "1001" when "101001101100",  -- brick
        "0101" when "101100111110",  -- block
        "0101" when "110000010000",  -- block
        "0010" when "110011100010",  -- death
        "1001" when "100011001001",  -- brick
        "1001" when "100110011011",  -- brick
        "1001" when "101001101101",  -- brick
        "0101" when "101100111111",  -- block
        "0101" when "110000010001",  -- block
        "0010" when "110011100011",  -- death
        "1001" when "011111111000",  -- brick
        "1001" when "100011001010",  -- brick
        "1001" when "100110011100",  -- brick
        "1001" when "101001101110",  -- brick
        "0101" when "101101000000",  -- block
        "0101" when "110000010010",  -- block
        "0010" when "110011100100",  -- death
        "1001" when "011111111001",  -- brick
        "1001" when "100011001011",  -- brick
        "1001" when "100110011101",  -- brick
        "1001" when "101001101111",  -- brick
        "0101" when "101101000001",  -- block
        "0101" when "110000010011",  -- block
        "0010" when "110011100101",  -- death
        "0010" when "110011100110",  -- death
        "0010" when "110011100111",  -- death
        "1001" when "011111111100",  -- brick
        "1001" when "100011001110",  -- brick
        "1001" when "100110100000",  -- brick
        "1001" when "101001110010",  -- brick
        "0101" when "101101000100",  -- block
        "0101" when "110000010110",  -- block
        "0010" when "110011101000",  -- death
        "1001" when "100011001111",  -- brick
        "1001" when "100110100001",  -- brick
        "1001" when "101001110011",  -- brick
        "0101" when "101101000101",  -- block
        "0101" when "110000010111",  -- block
        "0010" when "110011101001",  -- death
        "1001" when "100110100010",  -- brick
        "1001" when "101001110100",  -- brick
        "0101" when "101101000110",  -- block
        "0101" when "110000011000",  -- block
        "0010" when "110011101010",  -- death
        "1001" when "101001110101",  -- brick
        "0101" when "101101000111",  -- block
        "0101" when "110000011001",  -- block
        "0010" when "110011101011",  -- death
        "0101" when "101101001000",  -- block
        "0101" when "110000011010",  -- block
        "0010" when "110011101100",  -- death
        "0101" when "101101001001",  -- block
        "0101" when "110000011011",  -- block
        "0010" when "110011101101",  -- death
        "0101" when "101101001010",  -- block
        "0101" when "110000011100",  -- block
        "0010" when "110011101110",  -- death
        "0101" when "101101001011",  -- block
        "0101" when "110000011101",  -- block
        "0010" when "110011101111",  -- death
        "1001" when "100110101000",  -- brick
        "1001" when "101001111010",  -- brick
        "0101" when "101101001100",  -- block
        "0101" when "110000011110",  -- block
        "0010" when "110011110000",  -- death
        "1001" when "100110101001",  -- brick
        "1001" when "101001111011",  -- brick
        "0101" when "101101001101",  -- block
        "0101" when "110000011111",  -- block
        "0010" when "110011110001",  -- death
        "0101" when "101101001110",  -- block
        "0101" when "110000100000",  -- block
        "0010" when "110011110010",  -- death
        "0101" when "101101001111",  -- block
        "0101" when "110000100001",  -- block
        "0010" when "110011110011",  -- death
        "0101" when "101101010000",  -- block
        "0101" when "110000100010",  -- block
        "0010" when "110011110100",  -- death
        "1001" when "100000001001",  -- brick
        "0101" when "101101010001",  -- block
        "0101" when "110000100011",  -- block
        "0010" when "110011110101",  -- death
        -- all blocks except 'air' in screen 8 are below
        "1001" when "100000001010",  -- brick
        "0101" when "101101010010",  -- block
        "0101" when "110000100100",  -- block
        "0010" when "110011110110",  -- death
        "0101" when "100000001011",  -- block
        "0101" when "101101010011",  -- block
        "0101" when "110000100101",  -- block
        "0010" when "110011110111",  -- death
        "1001" when "100000001100",  -- brick
        "0101" when "101101010100",  -- block
        "0101" when "110000100110",  -- block
        "0010" when "110011111000",  -- death
        "0101" when "101101010101",  -- block
        "0101" when "110000100111",  -- block
        "0010" when "110011111001",  -- death
        "0101" when "101101010110",  -- block
        "0101" when "110000101000",  -- block
        "0010" when "110011111010",  -- death
        "0101" when "101101010111",  -- block
        "0101" when "110000101001",  -- block
        "0010" when "110011111011",  -- death
        "0101" when "101101011000",  -- block
        "0101" when "110000101010",  -- block
        "0010" when "110011111100",  -- death
        "1001" when "100110110101",  -- brick
        "1001" when "101010000111",  -- brick
        "0101" when "101101011001",  -- block
        "0101" when "110000101011",  -- block
        "0010" when "110011111101",  -- death
        "1001" when "100110110110",  -- brick
        "1001" when "101010001000",  -- brick
        "0101" when "101101011010",  -- block
        "0101" when "110000101100",  -- block
        "0010" when "110011111110",  -- death
        "0101" when "101101011011",  -- block
        "0101" when "110000101101",  -- block
        "0010" when "110011111111",  -- death
        "0101" when "101101011100",  -- block
        "0101" when "110000101110",  -- block
        "0010" when "110100000000",  -- death
        "0101" when "101101011101",  -- block
        "0101" when "110000101111",  -- block
        "0010" when "110100000001",  -- death
        "1001" when "101010001100",  -- brick
        "0101" when "101101011110",  -- block
        "0101" when "110000110000",  -- block
        "0010" when "110100000010",  -- death
        "1001" when "100110111011",  -- brick
        "1001" when "101010001101",  -- brick
        "0101" when "101101011111",  -- block
        "0101" when "110000110001",  -- block
        "0010" when "110100000011",  -- death
        "1001" when "100011101010",  -- brick
        "1001" when "100110111100",  -- brick
        "1001" when "101010001110",  -- brick
        "0101" when "101101100000",  -- block
        "0101" when "110000110010",  -- block
        "0010" when "110100000100",  -- death
        "1001" when "100000011001",  -- brick
        "1001" when "100011101011",  -- brick
        "1001" when "100110111101",  -- brick
        "1001" when "101010001111",  -- brick
        "0101" when "101101100001",  -- block
        "0101" when "110000110011",  -- block
        "0010" when "110100000101",  -- death
        "1001" when "011101001000",  -- brick
        "1001" when "100000011010",  -- brick
        "1001" when "100011101100",  -- brick
        "1001" when "100110111110",  -- brick
        "1001" when "101010010000",  -- brick
        "0101" when "101101100010",  -- block
        "0101" when "110000110100",  -- block
        "0010" when "110100000110",  -- death
        "1001" when "011001110111",  -- brick
        "1001" when "011101001001",  -- brick
        "1001" when "100000011011",  -- brick
        "1001" when "100011101101",  -- brick
        "1001" when "100110111111",  -- brick
        "1001" when "101010010001",  -- brick
        "0101" when "101101100011",  -- block
        "0101" when "110000110101",  -- block
        "0010" when "110100000111",  -- death
        "1001" when "010110100110",  -- brick
        "1001" when "011001111000",  -- brick
        "1001" when "011101001010",  -- brick
        "1001" when "100000011100",  -- brick
        "1001" when "100011101110",  -- brick
        "1001" when "100111000000",  -- brick
        "1001" when "101010010010",  -- brick
        "0101" when "101101100100",  -- block
        "0101" when "110000110110",  -- block
        "0010" when "110100001000",  -- death
        "1001" when "010011010101",  -- brick
        "1001" when "010110100111",  -- brick
        "1001" when "011001111001",  -- brick
        "1001" when "011101001011",  -- brick
        "1001" when "100000011101",  -- brick
        "1001" when "100011101111",  -- brick
        "1001" when "100111000001",  -- brick
        "1001" when "101010010011",  -- brick
        "0101" when "101101100101",  -- block
        "0101" when "110000110111",  -- block
        "0010" when "110100001001",  -- death
        "0101" when "101101100110",  -- block
        "0101" when "110000111000",  -- block
        "0010" when "110100001010",  -- death
        -- all blocks except 'air' in screen 9 are below
        "0101" when "101101100111",  -- block
        "0101" when "110000111001",  -- block
        "0010" when "110100001011",  -- death
        "0101" when "101101101000",  -- block
        "0101" when "110000111010",  -- block
        "0010" when "110100001100",  -- death
        "0101" when "101101101001",  -- block
        "0101" when "110000111011",  -- block
        "0010" when "110100001101",  -- death
        "0101" when "101101101010",  -- block
        "0101" when "110000111100",  -- block
        "0010" when "110100001110",  -- death
        "0101" when "101101101011",  -- block
        "0101" when "110000111101",  -- block
        "0010" when "110100001111",  -- death
        "0101" when "101101101100",  -- block
        "0101" when "110000111110",  -- block
        "0010" when "110100010000",  -- death
        "0101" when "101101101101",  -- block
        "0101" when "110000111111",  -- block
        "0010" when "110100010001",  -- death
        "0011" when "001001101000",  -- win
        "0011" when "001100111010",  -- win
        "0011" when "010000001100",  -- win
        "0011" when "010011011110",  -- win
        "0011" when "010110110000",  -- win
        "0011" when "011010000010",  -- win
        "0011" when "011101010100",  -- win
        "0011" when "100000100110",  -- win
        "0011" when "100011111000",  -- win
        "0011" when "100111001010",  -- win
        "1001" when "101010011100",  -- brick
        "0101" when "101101101110",  -- block
        "0101" when "110001000000",  -- block
        "0010" when "110100010010",  -- death
        "0101" when "101101101111",  -- block
        "0101" when "110001000001",  -- block
        "0010" when "110100010011",  -- death
        "0101" when "101101110000",  -- block
        "0101" when "110001000010",  -- block
        "0010" when "110100010100",  -- death
        "0101" when "101101110001",  -- block
        "0101" when "110001000011",  -- block
        "0010" when "110100010101",  -- death
        "0101" when "100000101010",  -- block
        "1001" when "100011111100",  -- brick
        "1001" when "100111001110",  -- brick
        "1001" when "101010100000",  -- brick
        "0101" when "101101110010",  -- block
        "0101" when "110001000100",  -- block
        "0010" when "110100010110",  -- death
        "0101" when "011010000111",  -- block
        "1001" when "011101011001",  -- brick
        "1001" when "100000101011",  -- brick
        "1001" when "100011111101",  -- brick
        "1001" when "100111001111",  -- brick
        "1001" when "101010100001",  -- brick
        "0101" when "101101110011",  -- block
        "0101" when "110001000101",  -- block
        "0010" when "110100010111",  -- death
        "0101" when "011101011010",  -- block
        "1001" when "100000101100",  -- brick
        "1001" when "100011111110",  -- brick
        "0101" when "100111010000",  -- block
        "0101" when "101010100010",  -- block
        "0101" when "101101110100",  -- block
        "0101" when "110001000110",  -- block
        "0010" when "110100011000",  -- death
        "0101" when "011010001001",  -- block
        "1001" when "011101011011",  -- brick
        "1001" when "100000101101",  -- brick
        "0101" when "100011111111",  -- block
        "0101" when "100111010001",  -- block
        "0101" when "101010100011",  -- block
        "0101" when "101101110101",  -- block
        "0101" when "110001000111",  -- block
        "0010" when "110100011001",  -- death
        "0101" when "011101011100",  -- block
        "1001" when "100000101110",  -- brick
        "1001" when "100100000000",  -- brick
        "0101" when "100111010010",  -- block
        "0101" when "101010100100",  -- block
        "0101" when "101101110110",  -- block
        "0101" when "110001001000",  -- block
        "0010" when "110100011010",  -- death
        "0101" when "011010001011",  -- block
        "1001" when "011101011101",  -- brick
        "1001" when "100000101111",  -- brick
        "1001" when "100100000001",  -- brick
        "1001" when "100111010011",  -- brick
        "1001" when "101010100101",  -- brick
        "0101" when "101101110111",  -- block
        "0101" when "110001001001",  -- block
        "0010" when "110100011011",  -- death
        "0101" when "100000110000",  -- block
        "1001" when "100100000010",  -- brick
        "1001" when "100111010100",  -- brick
        "1001" when "101010100110",  -- brick
        "0101" when "101101111000",  -- block
        "0101" when "110001001010",  -- block
        "0010" when "110100011100",  -- death
        "0101" when "101101111001",  -- block
        "0101" when "110001001011",  -- block
        "0010" when "110100011101",  -- death
        "0101" when "101101111010",  -- block
        "0101" when "110001001100",  -- block
        "0010" when "110100011110",  -- death
        "0101" when "101101111011",  -- block
        "0101" when "110001001101",  -- block
        "0010" when "110100011111",  -- death
        "0000" when others;  -- air

end lut;

