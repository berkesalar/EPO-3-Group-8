library ieee;
use ieee.std_logic_1164.all;
 
entity dabble is
    port (      A_in            : in std_logic_vector (3 downto 0);
                A_out           : out std_logic_vector (3 downto 0));
end dabble;