library ieee;
use ieee.std_logic_1164.all;

entity win_lut is
    port (
        addr    : in std_logic_vector(7 downto 0);
        blk_data: out std_logic
    );
end entity win_lut;

architecture lut of win_lut is

begin
    with addr select blk_data <= -- 0 = transparent/black, 1 = white
        '1' when "00000000",
        '0' when "00000001",
        '0' when "00000010",
        '0' when "00000011",
        '1' when "00000100",
        '0' when "00000101",
        '1' when "00000110",
        '1' when "00000111",
        '1' when "00001000",
        '0' when "00001001",
        '1' when "00001010",
        '0' when "00001011",
        '0' when "00001100",
        '1' when "00001101",
        '0' when "00001110",
        '1' when "00001111",
        '1' when "00010000",
        '1' when "00010001",
        '0' when "00010010",
        '0' when "00010011",
        '0' when "00010100",
        '1' when "00010101",
        '0' when "00010110",
        '0' when "00010111",
        '1' when "00011000",
        '0' when "00011001",
        '0' when "00011010",
        '1' when "00011011",
        '1' when "00011100",
        '0' when "00011101",
        '1' when "00011110",
        '0' when "00011111",
        '1' when "00100000",
        '1' when "00100001",
        '1' when "00100010",
        '0' when "00100011",
        '1' when "00100100",
        '0' when "00100101",
        '1' when "00100110",
        '0' when "00100111",
        '0' when "00101000",
        '1' when "00101001",
        '0' when "00101010",
        '0' when "00101011",
        '1' when "00101100",
        '0' when "00101101",
        '1' when "00101110",
        '1' when "00101111",
        '0' when "00110000",
        '1' when "00110001",
        '0' when "00110010",
        '1' when "00110011",
        '1' when "00110100",
        '0' when "00110101",
        '1' when "00110110",
        '1' when "00110111",
        '0' when "00111000",
        '0' when "00111001",
        '1' when "00111010",
        '0' when "00111011",
        '0' when "00111100",
        '1' when "00111101",
        '0' when "00111110",
        '0' when "00111111",
        '1' when "01000000",
        '0' when "01000001",
        '0' when "01000010",
        '0' when "01000011",
        '1' when "01000100",
        '0' when "01000101",
        '0' when "01000110",
        '0' when "01000111",
        '1' when "01001000",
        '0' when "01001001",
        '1' when "01001010",
        '1' when "01001011",
        '1' when "01001100",
        '0' when "01001101",
        '1' when "01001110",
        '0' when "01001111",
        '0' when "01010000",
        '1' when "01010001",
        '0' when "01010010",
        '1' when "01010011",
        '0' when "01010100",
        '0' when others;
end lut; 
