library ieee;
use ieee.std_logic_1164.all;

entity start_lut is
    port (
        addr    : in std_logic_vector(7 downto 0);
        blk_data: out std_logic
    );
end entity start_lut;

architecture lut of start_lut is

begin
    with addr select blk_data <= -- 0 = transparent/black, 1 = white
        '0' when "00000000",
        '1' when "00000001",
        '1' when "00000010",
        '1' when "00000011",
        '0' when "00000100",
        '1' when "00000101",
        '1' when "00000110",
        '1' when "00000111",
        '0' when "00001000",
        '0' when "00001001",
        '1' when "00001010",
        '1' when "00001011",
        '0' when "00001100",
        '0' when "00001101",
        '1' when "00001110",
        '1' when "00001111",
        '1' when "00010000",
        '0' when "00010001",
        '0' when "00010010",
        '1' when "00010011",
        '1' when "00010100",
        '1' when "00010101",
        '0' when "00010110",
        '0' when "00010111",
        '1' when "00011000",
        '1' when "00011001",
        '1' when "00011010",
        '0' when "00011011",
        '1' when "00011100",
        '0' when "00011101",
        '0' when "00011110",
        '0' when "00011111",
        '0' when "00100000",
        '0' when "00100001",
        '1' when "00100010",
        '0' when "00100011",
        '0' when "00100100",
        '1' when "00100101",
        '0' when "00100110",
        '0' when "00100111",
        '1' when "00101000",
        '0' when "00101001",
        '1' when "00101010",
        '0' when "00101011",
        '0' when "00101100",
        '1' when "00101101",
        '0' when "00101110",
        '0' when "00101111",
        '1' when "00110000",
        '0' when "00110001",
        '0' when "00110010",
        '1' when "00110011",
        '0' when "00110100",
        '0' when "00110101",
        '0' when "00110110",
        '1' when "00110111",
        '1' when "00111000",
        '1' when "00111001",
        '1' when "00111010",
        '1' when "00111011",
        '0' when "00111100",
        '0' when "00111101",
        '1' when "00111110",
        '0' when "00111111",
        '0' when "01000000",
        '1' when "01000001",
        '1' when "01000010",
        '1' when "01000011",
        '1' when "01000100",
        '0' when "01000101",
        '1' when "01000110",
        '0' when "01000111",
        '1' when "01001000",
        '1' when "01001001",
        '0' when "01001010",
        '0' when "01001011",
        '1' when "01001100",
        '0' when "01001101",
        '0' when "01001110",
        '0' when "01001111",
        '0' when "01010000",
        '1' when "01010001",
        '1' when "01010010",
        '0' when "01010011",
        '0' when "01010100",
        '0' when "01010101",
        '0' when "01010110",
        '1' when "01010111",
        '0' when "01011000",
        '0' when "01011001",
        '1' when "01011010",
        '0' when "01011011",
        '0' when "01011100",
        '1' when "01011101",
        '0' when "01011110",
        '0' when "01011111",
        '1' when "01100000",
        '0' when "01100001",
        '1' when "01100010",
        '1' when "01100011",
        '0' when "01100100",
        '0' when "01100101",
        '0' when "01100110",
        '0' when "01100111",
        '1' when "01101000",
        '0' when "01101001",
        '0' when "01101010",
        '0' when "01101011",
        '0' when "01101100",
        '0' when "01101101",
        '0' when "01101110",
        '0' when "01101111",
        '1' when "01110000",
        '1' when "01110001",
        '1' when "01110010",
        '0' when "01110011",
        '0' when "01110100",
        '0' when "01110101",
        '1' when "01110110",
        '0' when "01110111",
        '0' when "01111000",
        '1' when "01111001",
        '0' when "01111010",
        '0' when "01111011",
        '1' when "01111100",
        '0' when "01111101",
        '1' when "01111110",
        '0' when "01111111",
        '1' when "10000000",
        '1' when "10000001",
        '0' when "10000010",
        '0' when "10000011",
        '1' when "10000100",
        '0' when "10000101",
        '0' when "10000110",
        '0' when "10000111",
        '0' when "10001000",
        '1' when "10001001",
        '0' when "10001010",
        '0' when "10001011",
        '0' when others;
        
end lut; 
