library ieee;
use ieee.std_logic_1164.all;

entity game_over_lut is
    port (
        addr    : in std_logic_vector(7 downto 0);
        blk_data: out std_logic
    );
end entity game_over_lut;

architecture lut of game_over_lut is

begin
    with addr select blk_data <= -- 0 = transparent/black, 1 = white
        '0' when "00000000",
        '1' when "00000001",
        '1' when "00000010",
        '1' when "00000011",
        '0' when "00000100",
        '0' when "00000101",
        '1' when "00000110",
        '1' when "00000111",
        '0' when "00001000",
        '0' when "00001001",
        '1' when "00001010",
        '0' when "00001011",
        '0' when "00001100",
        '0' when "00001101",
        '1' when "00001110",
        '0' when "00001111",
        '1' when "00010000",
        '1' when "00010001",
        '1' when "00010010",
        '1' when "00010011",
        '0' when "00010100",
        '0' when "00010101",
        '0' when "00010110",
        '0' when "00010111",
        '1' when "00011000",
        '1' when "00011001",
        '0' when "00011010",
        '0' when "00011011",
        '1' when "00011100",
        '0' when "00011101",
        '0' when "00011110",
        '0' when "00011111",
        '1' when "00100000",
        '0' when "00100001",
        '1' when "00100010",
        '1' when "00100011",
        '1' when "00100100",
        '1' when "00100101",
        '0' when "00100110",
        '1' when "00100111",
        '1' when "00101000",
        '1' when "00101001",
        '0' when "00101010",
        '0' when "00101011",
        '1' when "00101100",
        '1' when "00101101",
        '1' when "00101110",
        '0' when "00101111",
        '0' when "00110000",
        '0' when "00110001",
        '0' when "00110010",
        '1' when "00110011",
        '0' when "00110100",
        '0' when "00110101",
        '1' when "00110110",
        '0' when "00110111",
        '1' when "00111000",
        '1' when "00111001",
        '0' when "00111010",
        '1' when "00111011",
        '1' when "00111100",
        '0' when "00111101",
        '1' when "00111110",
        '0' when "00111111",
        '0' when "01000000",
        '0' when "01000001",
        '0' when "01000010",
        '0' when "01000011",
        '0' when "01000100",
        '1' when "01000101",
        '0' when "01000110",
        '0' when "01000111",
        '1' when "01001000",
        '0' when "01001001",
        '1' when "01001010",
        '0' when "01001011",
        '0' when "01001100",
        '0' when "01001101",
        '1' when "01001110",
        '0' when "01001111",
        '1' when "01010000",
        '0' when "01010001",
        '0' when "01010010",
        '0' when "01010011",
        '0' when "01010100",
        '1' when "01010101",
        '0' when "01010110",
        '0' when "01010111",
        '1' when "01011000",
        '0' when "01011001",
        '1' when "01011010",
        '1' when "01011011",
        '1' when "01011100",
        '0' when "01011101",
        '1' when "01011110",
        '1' when "01011111",
        '0' when "01100000",
        '1' when "01100001",
        '1' when "01100010",
        '1' when "01100011",
        '1' when "01100100",
        '0' when "01100101",
        '1' when "01100110",
        '0' when "01100111",
        '1' when "01101000",
        '0' when "01101001",
        '1' when "01101010",
        '0' when "01101011",
        '1' when "01101100",
        '1' when "01101101",
        '1' when "01101110",
        '0' when "01101111",
        '0' when "01110000",
        '0' when "01110001",
        '0' when "01110010",
        '1' when "01110011",
        '0' when "01110100",
        '0' when "01110101",
        '1' when "01110110",
        '0' when "01110111",
        '1' when "01111000",
        '0' when "01111001",
        '0' when "01111010",
        '0' when "01111011",
        '1' when "01111100",
        '0' when "01111101",
        '1' when "01111110",
        '1' when "01111111",
        '1' when "10000000",
        '0' when "10000001",
        '0' when "10000010",
        '1' when "10000011",
        '0' when "10000100",
        '1' when "10000101",
        '1' when "10000110",
        '0' when "10000111",
        '1' when "10001000",
        '0' when "10001001",
        '1' when "10001010",
        '0' when "10001011",
        '0' when "10001100",
        '1' when "10001101",
        '0' when "10001110",
        '1' when "10001111",
        '0' when "10010000",
        '0' when "10010001",
        '1' when "10010010",
        '0' when "10010011",
        '1' when "10010100",
        '0' when "10010101",
        '0' when "10010110",
        '0' when "10010111",
        '1' when "10011000",
        '0' when "10011001",
        '1' when "10011010",
        '0' when "10011011",
        '0' when "10011100",
        '0' when "10011101",
        '0' when "10011110",
        '0' when "10011111",
        '0' when "10100000",
        '1' when "10100001",
        '0' when "10100010",
        '0' when "10100011",
        '1' when "10100100",
        '0' when "10100101",
        '0' when "10100110",
        '1' when "10100111",
        '0' when "10101000",
        '1' when "10101001",
        '0' when "10101010",
        '0' when "10101011",
        '1' when "10101100",
        '0' when "10101101",
        '0' when "10101110",
        '0' when "10101111",
        '0' when "10110000",
        '1' when "10110001",
        '1' when "10110010",
        '0' when "10110011",
        '0' when "10110100",
        '0' when "10110101",
        '0' when "10110110",
        '0' when "10110111",
        '0' when "10111000",
        '1' when "10111001",
        '1' when "10111010",
        '1' when "10111011",
        '0' when "10111100",
        '1' when "10111101",
        '0' when "10111110",
        '0' when "10111111",
        '1' when "11000000",
        '0' when "11000001",
        '1' when "11000010",
        '0' when "11000011",
        '0' when "11000100",
        '0' when "11000101",
        '1' when "11000110",
        '0' when "11000111",
        '1' when "11001000",
        '1' when "11001001",
        '1' when "11001010",
        '1' when "11001011",
        '0' when "11001100",
        '0' when "11001101",
        '0' when "11001110",
        '0' when "11001111",
        '1' when "11010000",
        '1' when "11010001",
        '0' when "11010010",
        '0' when "11010011",
        '0' when "11010100",
        '0' when "11010101",
        '1' when "11010110",
        '0' when "11010111",
        '0' when "11011000",
        '0' when "11011001",
        '1' when "11011010",
        '1' when "11011011",
        '1' when "11011100",
        '1' when "11011101",
        '0' when "11011110",
        '1' when "11011111",
        '0' when "11100000",
        '1' when "11100001",
        '1' when "11100010",
        '0' when "11100011",
        '1' when "11100100",
        '0' when "11100101",
        '0' when others;
    
end lut; 
